*Four pixel digital camera

.param proc_delta = 1.0
.param vt_shift = 0.0

* p18 model card
.MODEL NMOS NMOS  								
+ VERSION	=	3.1						
+ LEVEL	=	49	NOIMOD	=	1	TNOM	=	2.70E+01
+ TOX	=	'4.1E-9/proc_delta'	XJ	=	1.00E-07	NCH	=	2.33E+17
+ VTH0	=	'0.36+vt_shift'	K1	=	5.84E-01	K2	=	4.14E-03
+ K3	=	1.01E-03	K3B	=	2.20E+00	W0	=	1.00E-07
+ NLX	=	1.81E-07	DVT0W	=	0.00E+00	DVT1W	=	0.00E+00
+ DVT2W	=	0.00E+00	DVT0	=	1.73E+00	DVT1	=	4.38E-01
+ DVT2	=	-3.70E-04	U0	=	'260*proc_delta*proc_delta'	UA	=	-1.38E-09
+ UB	=	2.26E-18	UC	=	5.46E-11	VSAT	=	1.03E+05
+ A0	=	1.92E+00	AGS	=	4.20E-01	B0	=	-1.52E-09
+ B1	=	-9.92E-08	KETA	=	-7.16E-03	A1	=	6.61E-04
+ A2	=	8.89E-01	RDSW	=	1.12E+02	PRWG	=	4.92E-01
+ PRWB	=	-2.02E-01	WR	=	1.00E+00	WINT	=	7.12E-09
+ LINT	=	1.12E-08	XL	=	-2.00E-08	XW	=	-1.00E-08
+ DWG	=	-3.82E-09	DWB	=	8.63E-09	VOFF	=	-8.82E-02
+ NFACTOR	=	2.30E+00	CIT	=	0.00E+00	CDSC	=	2.40E-04
+ CDSCD	=	0.00E+00	CDSCB	=	0.00E+00	ETA0	=	3.13E-03
+ ETAB	=	1.00E+00	DSUB	=	2.25E-02	PCLM	=	7.20E-01
+ PDIBLC1	=	2.15E-01	PDIBLC2	=	2.23E-03	PDIBLCB	=	1.00E-01
+ DROUT	=	8.01E-01	PSCBE1	=	5.44E+08	PSCBE2	=	1.00E-03
+ PVAG	=	1.00E-12	DELTA	=	1.00E-02	RSH	=	6.78E+00
+ MOBMOD	=	1.00E+00	PRT	=	0.00E+00	UTE	=	-1.50E+00
+ KT1	=	-1.10E-01	KT1L	=	0.00E+00	KT2	=	2.19E-02
+ UA1	=	4.28E-09	UB1	=	-7.62E-18	UC1	=	-5.57E-11
+ AT	=	3.30E+04	WL	=	0.00E+00	WLN	=	1.00E+00
+ WW	=	0.00E+00	WWN	=	1.00E+00	WWL	=	0.00E+00
+ LL	=	0.00E+00	LLN	=	1.00E+00	LW	=	0.00E+00
+ LWN	=	1.00E+00	LWL	=	0.00E+00	CAPMOD	=	2.00E+00
+ XPART	=	5.00E-01	CGDO	=	6.98E-10	CGSO	=	7.03E-10
+ CGBO	=	1.00E-12	CJ	=	'9.8e-4/proc_delta'	PB	=	7.34E-01
+ MJ	=	3.63E-01	CJSW	=	'2.4e-10/proc_delta'	PBSW	=	4.71E-01
+ MJSW	=	1.00E-01	CJSWG	=	3.29E-10	PBSWG	=	4.66E-01
+ MJSWG	=	1.00E-01	CF	=	0.00E+00	PVTH0	=	-7.16E-04
+ PRDSW	=	-6.66E-01	PK2	=	5.92E-04	WKETA	=	2.14E-04
+ LKETA	=	-1.51E-02	PU0	=	3.36E+00	PUA	=	-1.31E-11
+ PUB	=	0.00E+00	PVSAT	=	1.25E+03	PETA0	=	1.00E-04
+ PKETA	=	6.45E-04	KF	=	4.46E-29			

.MODEL PMOS PMOS  								
+ VERSION	=	3.1						
+ LEVEL	=	49	NOIMOD	=	1			
+ TNOM	=	2.70E+01	TOX	=	'4.1E-9/proc_delta'	XJ	=	1.00E-07
+ NCH	=	4.12E+17	VTH0	=	'-0.39-vt_shift'	K1	=	5.50E-01
+ K2	=	3.50E-02	K3	=	0.00E+00	K3B	=	1.20E+01
+ W0	=	1.00E-06	NLX	=	1.25E-07	DVT0W	=	0.00E+00
+ DVT1W	=	0.00E+00	DVT2W	=	0.00E+00	DVT0	=	5.53E-01
+ DVT1	=	2.46E-01	DVT2	=	1.00E-01	U0	=	'110*proc_delta*proc_delta'
+ UA	=	1.44E-09	UB	=	2.29E-21	UC	=	-1.00E-10
+ VSAT	=	1.95E+05	A0	=	1.72E+00	AGS	=	3.80E-01
+ B0	=	5.87E-07	B1	=	1.44E-06	KETA	=	2.21E-02
+ A1	=	4.66E-01	A2	=	3.00E-01	RDSW	=	3.11E+02
+ PRWG	=	5.00E-01	PRWB	=	1.64E-02	WR	=	1.00E+00
+ WINT	=	0.00E+00	LINT	=	2.00E-08	XL	=	-2.00E-08
+ XW	=	-1.00E-08	DWG	=	-3.49E-08	DWB	=	1.22E-09
+ VOFF	=	-9.80E-02	NFACTOR	=	2.00E+00	CIT	=	0.00E+00
+ CDSC	=	2.40E-04	CDSCD	=	0.00E+00	CDSCB	=	0.00E+00
+ ETA0	=	1.12E-03	ETAB	=	-4.79E-04	DSUB	=	1.60E-03
+ PCLM	=	1.50E+00	PDIBLC1	=	3.00E-02	PDIBLC2	=	-1.01E-05
+ PDIBLCB	=	1.00E-01	DROUT	=	1.56E-03	PSCBE1	=	4.91E+09
+ PSCBE2	=	1.64E-09	PVAG	=	3.48E+00	DELTA	=	1.00E-02
+ RSH	=	7.69E+00	MOBMOD	=	1.00E+00	PRT	=	0.00E+00
+ UTE	=	-1.49E+00	KT1	=	-1.09E-01	KT1L	=	0.00E+00
+ KT2	=	2.18E-02	UA1	=	4.27E-09	UB1	=	-7.68E-18
+ UC1	=	-5.57E-11	AT	=	3.31E+04	WL	=	0.00E+00
+ WLN	=	1.00E+00	WW	=	0.00E+00	WWN	=	1.00E+00
+ WWL	=	0.00E+00	LL	=	0.00E+00	LLN	=	1.00E+00
+ LW	=	0.00E+00	LWN	=	1.00E+00	LWL	=	0.00E+00
+ CAPMOD	=	2.00E+00	XPART	=	5.00E-01	CGDO	=	6.88E-10
+ CGSO	=	6.85E-10	CGBO	=	1.00E-12	CJ	=	'1.2e-3/proc_delta'
+ PB	=	8.70E-01	MJ	=	4.20E-01	CJSW	=	'2.4e-10/proc_delta'
+ PBSW	=	8.00E-01	MJSW	=	3.57E-01	CJSWG	=	4.24E-10
+ PBSWG	=	8.00E-01	MJSWG	=	3.56E-01	CF	=	0.00E+00
+ PVTH0	=	3.53E-03	PRDSW	=	1.02E+01	PK2	=	3.35E-03
+ WKETA	=	3.52E-02	LKETA	=	-2.06E-03	PU0	=	-2.19E+00
+ PUA	=	-7.63E-11	PUB	=	9.91E-22	PVSAT	=	5.00E+01
+ PKETA	=	-6.41E-03	KF	=	1.29E-29	PETA0	=	7.31E-05


.param Ipd_1 = 50p
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 30m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

.param minW=1.08u
.param maxW=5.04u
.param maxL=1.08u
.param minL=0.36u

.param MswitchW=minW
.param MswitchL=maxL
.param MbufferW=maxW
.param MbufferL=minL

.param MactiveLoadW=minW
.param MactiveLoadL=maxL
.param CC_cap=3p

.param CS_cap=2p

.subckt PhotoDiode  VDD N1_R1C1 
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1            ! Photo current source
d1 N1_R1C1 VDD dwell 1                        ! Reverse biased Diode
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40 ! Diode model
Cd1 N1_R1C1 VDD 30f                           ! Photo diode capacitor
.ends

.subckt pixel VDD VSS EXPOSE ERASE NRE OUT N2
xPhotoDiode VDD 1 PhotoDiode

M1 1 EXPOSE N2 VSS NMOS W=MswitchW L=MswitchL
M2 N2 ERASE VSS VSS NMOS W=MswitchW L=MswitchL

CS N2 VSS CS_cap

M3 3 N2 VSS VDD PMOS W=MbufferW L=MbufferL
M4 OUT NRE 3 VDD PMOS W=MswitchW L=MswitchL
.ends

.subckt load VDD VSS OUT
MC VDD OUT OUT VDD PMOS W=MactiveLoadW L=MactiveLoadL
CC OUT VSS CC_cap
.ends

xPixel_11 1 0 2 3 4 6  8 pixel
xPixel_12 1 0 2 3 4 7  9 pixel
xPixel_21 1 0 2 3 5 6 10 pixel
xPixel_22 1 0 2 3 5 7 11 pixel

xLoad1 1 0 6 load
xLoad2 1 0 7 load

VDD 1 0 dc VDD

vEXPOSE 2 0 dc 0 pulse(0v VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
vERASE  3 0 dc 0 pulse(0v VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)

vNRE1 4 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
vNRE2 5 0 dc 0 pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

*.plot TRAN V(6)
*.plot TRAN V(7)
.plot TRAN V(2) V(3) V(4) V(5) V(6) V(8)
*.plot TRAN V(4) V(5)
*.plot TRAN V(8)

.tran 20n 20m